module imm_gen (
    input [31:0] instruction,
    input [2:0] imm_sel,
    output reg [31:0] immediate
);

    localparam IMM_I = 3'b000;
    localparam IMM_S = 3'b001;
    localparam IMM_B = 3'b010;
    localparam IMM_U = 3'b011;
    localparam IMM_J = 3'b100;

    always @(*) begin
        case (imm_sel)
            IMM_I: immediate = {{20{instruction[31]}}, instruction[31:20]};

            IMM_S: immediate = {{20{instruction[31]}}, instruction[31:25], instruction[11:7]};

            IMM_B: immediate = {{19{instruction[31]}}, instruction[31], instruction[7],
                               instruction[30:25], instruction[11:8], 1'b0};

            IMM_U: immediate = {instruction[31:12], 12'b0};

            IMM_J: immediate = {{11{instruction[31]}}, instruction[31], instruction[19:12],
                               instruction[20], instruction[30:21], 1'b0};

            default: immediate = 32'd0;
        endcase
    end

endmodule
